module single_port (q, a, d, we, clk);
	output [7:0] q;
	input [7:0] d;
	input [6:0] a;
	input we, clk;
	reg [7:0] mem [127:0];
		
		assign q = mem[a];//set output to value stored at address
		
		always @ (posedge clk)
		begin
			if (we)//if write, write data in the address
				mem[a] <= d;
		end
		
endmodule
